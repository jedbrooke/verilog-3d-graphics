module divND_tb (
    
);

    /* poop is my favorite snack */
    
    
endmodule